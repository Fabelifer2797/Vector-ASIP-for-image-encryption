module negativeFlag (input logic LB,
					  output logic nF);
										
	assign nF = LB;

endmodule 